
module forward #(
  parameter [31:0] W = 16,
  parameter [31:0] N = 2,
  parameter [31:0] Q = 8
)(
  input clk,
  input rst,
  // Input connection slaves
  input [N-1:0] s_i_stb,
  input [N*W-1:0] s_i_dat,
  output [N-1:0] s_i_rdy,
  // Output connection master
  input m_o_rdy,
  output m_o_stb,
  output [W-1:0] m_o_dat,
  // Memory data slave
  input s_d_stb,
  input [W-1:0] s_d_dat,
  output s_d_rdy,
  // Memory address master
  input m_a_rdy,
  output m_a_stb,
  output [$clog2(N)-1:0] m_a_dat
);
  wire mux_stb;
  wire mux_rdy;
  wire [$clog2(N)+W-1:0] mux_dat;

  wire sep_stb;
  wire sep_rdy;
  wire [W-1:0] sep_dat;

  wire cmb_stb;
  wire cmb_rdy;
  wire [2*W-1:0] cmb_dat;

  wire mul_stb;
  wire mul_rdy;
  wire [2*W-1:0] mul_dat;

  wire acc_stb;
  wire acc_rdy;
  wire [2*W-1:0] acc_dat;

  wire [2*W-1:0] sat_dat;

  wire [W-$clog2(N):0] nc;
  wire unused = &{1'b0,
    nc,
    sat_dat[W+:W],
  1'b0};

  multiplex #(W, N) mux (
    .s_stb(s_i_stb),
    .s_dat(s_i_dat),
    .s_rdy(s_i_rdy),
    .m_rdy(mux_rdy),
    .m_stb(mux_stb),
    .m_dat(mux_dat)
  );

  seperate #(W) sep (
    .clk(clk),
    .rst(rst),
    .s_stb(mux_stb),
    .s_dat({{(W-$clog2(N)){1'bx}}, mux_dat}),
    .s_rdy(mux_rdy),
    .m_rdy({m_a_rdy, sep_rdy}),
    .m_stb({m_a_stb, sep_stb}),
    .m_dat({nc[1+:W-$clog2(N)], m_a_dat, sep_dat})
  );

  combine #(W) cmb (
    .s_stb({s_d_stb, sep_stb}),
    .s_dat({s_d_dat, sep_dat}),
    .s_rdy({s_d_rdy, sep_rdy}),
    .m_rdy(cmb_rdy),
    .m_stb(cmb_stb),
    .m_dat(cmb_dat)
  );

  multiply #(W, Q) mul (
    .clk(clk),
    .rst(rst),
    .s_stb(cmb_stb),
    .s_dat(cmb_dat),
    .s_rdy(cmb_rdy),
    .m_rdy(mul_rdy),
    .m_stb(mul_stb),
    .m_dat(mul_dat)
  );

  accumulate #(2*W) acc (
    .clk(clk),
    .rst(rst),
    .s_stb(mul_stb),
    .s_dat(mul_dat),
    .s_rdy(mul_rdy),
    .m_rdy(acc_rdy),
    .m_stb(acc_stb),
    .m_dat(acc_dat)
  );

  saturate #(2*W, W) sat (acc_dat, sat_dat);

  decimate #(W, N+1) dec (
    .clk(clk),
    .rst(rst),
    .s_stb(acc_stb),
    .s_dat(sat_dat[0+:W]),
    .s_rdy(acc_rdy),
    .m_rdy(m_o_rdy),
    .m_stb(m_o_stb),
    .m_dat(m_o_dat)
  );

endmodule
